`timescale 1ns / 1ps

module ControlALU(
    );


endmodule
