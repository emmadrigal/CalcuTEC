`timescale 1ns / 1ps

module PC_register(
    );


endmodule
