`timescale 1ns / 1ps

module ARMProcessor(
    );
	 
	 



endmodule
