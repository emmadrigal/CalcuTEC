`timescale 1ns / 1ps

module Mux2x1(
    );


endmodule
