`timescale 1ns / 1ps

module assemblytest;

	// Inputs
	reg clk;
	reg [31:0] datoA;
	reg [31:0] datoB;
	reg [2:0] operacion;
	reg start;

	// Outputs
	wire [31:0] resultado;
	wire ready;
	wire error;

	// Instantiate the Unit Under Test (UUT)
	Ensamblador uut (
		.clk(clk),
		.datoA(datoA), 
		.datoB(datoB), 
		.operacion(operacion), 
		.start(start), 
		.resultado(resultado), 
		.ready(ready), 
		.error(error)
	);

	initial begin
		// Initialize Inputs
		datoA = 0;
		datoB = 0;
		operacion = 0;
		start = 0;
		clk = 0;

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here
		#10; datoA = 5; datoB = 500; operacion = 4; start = 0;
		#10; start = 1; 
		#5; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;
		#1; clk = 1;
		#1; clk = 0;


	end
      
endmodule

