`timescale 1ns / 1ps

module TOP(
    );



endmodule
